

entity radio is
    port(
        [I/Os]
    );
end entity radio;