entity top_red is

end entity top_red;